library verilog;
use verilog.vl_types.all;
entity TB_CPU is
end TB_CPU;
